module ALU(
